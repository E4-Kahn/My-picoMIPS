`define LD   3'b000
`define BNE  3'b001
`define BEQ  3'b010
`define ADD  3'b100
`define ADDI 3'b101
`define MUL  3'b110
`define RLD   3'b000
`define RADD  3'b100
`define RADDI 3'b101
`define RMUL  3'b110
`define RBEQ  3'b010
`define RBNE  3'b001